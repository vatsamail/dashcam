package dashcam_uvm_agents_pkg;
  // Wishbone agent placeholder.
endpackage
