package dashcam_uvm_env_pkg;
  // UVM environment placeholder for Questa/Xcelium integration.
endpackage
