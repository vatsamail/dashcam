package dashcam_uvm_seq_pkg;
  // UVM sequence library placeholder.
endpackage
