package dashcam_uvm_tests_pkg;
  // UVM smoke test placeholder.
endpackage
